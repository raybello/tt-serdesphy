
interface sys_if;
    logic clk, rst_n;
    logic [31:0] pins;

endinterface
