/*
 * SerDes PHY Physical Medium Attachment
 * The PMA receives and transmits high-speed serial data on the serial lanes
 * Integrates PLL, CDR, Serializer, Deserializer, and differential I/O
 */

module serdesphy_pma(
    // Clock and Reset
    input  wire       clk_ref_24m,        // 24 MHz reference clock
    input  wire       rst_n,              // Global reset (active-low)
    input  wire       clk_240m_tx,        // 240 MHz TX clock (from outside, for compat)
    input  wire       clk_240m_rx,        // 240 MHz RX clock (from outside, for compat)

    // Power Control
    input  wire       analog_iso_n,       // Analog isolation (active-low)
    input  wire       analog_reset_n,     // Analog reset (active-low)

    // PLL Interface
    input  wire       pll_enable,         // PLL enable
    input  wire       pll_reset_n,        // PLL reset (active-low)
    input  wire       pll_bypass_en,      // PLL bypass enable
    input  wire [3:0] pll_vco_trim,       // PLL VCO trim
    input  wire [1:0] pll_cp_current,     // PLL charge pump current
    input  wire       pll_iso_n,          // PLL isolation (active-low)

    // PLL Status
    output wire       pll_lock_raw,       // Raw PLL lock
    output wire       pll_vco_ok,         // VCO OK indication
    output wire       pll_cp_ok,          // Charge pump OK indication

    // Clock Outputs (generated by PMA)
    output wire       clk_240m_pll,       // 240 MHz clock from PLL
    output wire       clk_240m_cdr,       // 240 MHz clock from CDR

    // TX Serializer Interface
    input  wire       serializer_enable,  // Serializer enable
    input  wire       serializer_clock,   // Serializer clock
    input  wire       serializer_reset_n, // Serializer reset (active-low)
    input  wire       serializer_data,    // Data to serializer
    input  wire       serializer_bypass,  // Serializer bypass (test mode)

    // Serializer Status
    output wire       serializer_ready,   // Serializer ready flag
    output wire       serializer_error,   // Serializer error flag
    output wire       serializer_active,  // Serializer active status
    output wire       serializer_status,  // Serializer status

    // RX Deserializer Interface
    input  wire       deserializer_enable,// Deserializer enable
    input  wire       deserializer_clock, // Deserializer clock reference
    input  wire       deserializer_reset_n,// Deserializer reset (active-low)
    input  wire       deserializer_bypass,// Deserializer bypass (test mode)

    // CDR Control
    input  wire [2:0] cdr_gain,           // CDR loop gain
    input  wire       cdr_fast_lock,      // CDR fast lock enable
    input  wire       cdr_rst,            // CDR reset

    // Deserializer Status
    output wire       deserializer_ready, // Deserializer ready flag
    output wire       deserializer_lock,  // Deserializer lock status (CDR lock)
    output wire       deserializer_error, // Deserializer error flag
    output wire       deserializer_active,// Deserializer active status
    output wire       deserializer_status,// Deserializer status
    output wire       deserializer_data,  // Serial data from deserializer

    // Differential TX Outputs
    output wire       txp,                // TX positive differential output
    output wire       txn,                // TX negative differential output

    // Differential RX Inputs
    input  wire       rxp,                // RX positive differential input
    input  wire       rxn,                // RX negative differential input

    // Loopback Control
    input  wire       lpbk_en,            // Loopback enable

    // Debug Interface
    input  wire       dbg_ana             // Debug analog control
);

    // =========================================================================
    // Internal Signals
    // =========================================================================

    wire analog_en;
    assign analog_en = analog_iso_n && analog_reset_n;

    // PLL signals
    wire       pll_clk_240m;
    wire [7:0] pll_vco_control;

    // TX path signals
    wire       tx_serial_out;
    wire       tx_driver_txp, tx_driver_txn;
    wire       serializer_busy;
    wire       serializer_data_ready;

    // Loopback signals
    wire       lpbk_rxp, lpbk_rxn;

    // RX path signals
    wire       rx_serial_data;
    wire       rx_signal_detected;
    wire [7:0] cdr_vco_control;
    wire       cdr_lock_int;
    wire       cdr_clk_240m;
    wire       cdr_vco_ready;
    wire [15:0] deser_parallel_out;
    wire       deser_data_valid;
    wire       deser_busy;

    // =========================================================================
    // PLL - Generates 240 MHz TX clock
    // =========================================================================

    serdesphy_ana_pll u_pll (
        .clk_ref_24m    (clk_ref_24m),
        .rst_n          (rst_n && analog_reset_n),
        .pll_rst        (!pll_reset_n),
        .pll_bypass     (pll_bypass_en),
        .enable         (pll_enable && analog_en),
        .vco_trim       (pll_vco_trim),
        .cp_current     (pll_cp_current),
        .clk_240m_out   (pll_clk_240m),
        .pll_lock       (pll_lock_raw),
        .vco_control    (pll_vco_control)
    );

    // PLL status
    assign pll_vco_ok = pll_lock_raw;  // VCO OK when PLL locked
    assign pll_cp_ok = pll_enable && analog_en;  // CP OK when enabled
    assign clk_240m_pll = pll_clk_240m;

    // =========================================================================
    // TX Path - Serializer and Differential Driver
    // =========================================================================

    // For now, use direct serial data pass-through since TX top handles serialization
    // The analog serializer is for future use with parallel data interface

    // TX Differential Driver
    serdesphy_ana_tx_differential_driver u_tx_driver (
        .clk            (pll_clk_240m),
        .rst_n          (rst_n && analog_reset_n && serializer_reset_n),
        .enable         (serializer_enable && analog_en),
        .serial_data    (serializer_data),
        .iso_en         (!analog_iso_n),
        .lpbk_en        (lpbk_en),
        .txp            (tx_driver_txp),
        .txn            (tx_driver_txn)
    );

    // Serializer status - simplified for direct serial mode
    assign serializer_ready = serializer_enable && analog_en && pll_lock_raw;
    assign serializer_error = 1'b0;
    assign serializer_active = serializer_enable && analog_en;
    assign serializer_status = serializer_ready;

    // TX outputs
    assign txp = tx_driver_txp;
    assign txn = tx_driver_txn;

    // =========================================================================
    // Loopback Switch
    // =========================================================================

    serdesphy_ana_loopback_switch u_loopback (
        .clk            (pll_clk_240m),
        .rst_n          (rst_n && analog_reset_n),
        .enable         (analog_en),
        .lpbk_en        (lpbk_en),
        .txp            (tx_driver_txp),
        .txn            (tx_driver_txn),
        .lpbk_rxp       (lpbk_rxp),
        .lpbk_rxn       (lpbk_rxn)
    );

    // =========================================================================
    // RX Path - Differential Receiver, CDR, and Deserializer
    // =========================================================================

    // RX Differential Receiver
    serdesphy_ana_rx_differential_receiver u_rx_receiver (
        .clk            (cdr_clk_240m),
        .rst_n          (rst_n && analog_reset_n && deserializer_reset_n),
        .enable         (deserializer_enable && analog_en),
        .rxp            (rxp),
        .rxn            (rxn),
        .iso_en         (!analog_iso_n),
        .lpbk_en        (lpbk_en),
        .lpbk_txp       (lpbk_rxp),
        .lpbk_txn       (lpbk_rxn),
        .serial_data    (rx_serial_data),
        .signal_detected(rx_signal_detected)
    );

    // CDR - Clock Data Recovery
    serdesphy_ana_cdr u_cdr (
        .clk_240m_rx    (cdr_clk_240m),
        .rst_n          (rst_n && analog_reset_n),
        .cdr_rst        (cdr_rst),
        .enable         (deserializer_enable && analog_en),
        .cdr_gain       (cdr_gain),
        .cdr_fast_lock  (cdr_fast_lock),
        .serial_data    (rx_serial_data),
        .vco_control    (cdr_vco_control),
        .cdr_lock       (cdr_lock_int),
        .phase_detector ()  // Not connected - internal debug
    );

    // CDR VCO - Generates recovered clock
    serdesphy_ana_cdr_vco u_cdr_vco (
        .rst_n          (rst_n && analog_reset_n),
        .enable         (deserializer_enable && analog_en),
        .cdr_control    (cdr_vco_control),
        .vco_out        (cdr_clk_240m),
        .vco_ready      (cdr_vco_ready)
    );

    assign clk_240m_cdr = cdr_clk_240m;

    // Deserializer status
    assign deserializer_ready = deserializer_enable && analog_en && cdr_vco_ready;
    assign deserializer_lock = cdr_lock_int;
    assign deserializer_error = 1'b0;
    assign deserializer_active = deserializer_enable && analog_en && rx_signal_detected;
    assign deserializer_status = cdr_lock_int;
    assign deserializer_data = rx_serial_data;

endmodule